//-------------------------------------------------------------------------
 //DUT+testbench+assertion
//-----------------------------------------------------------------------------------------------------------------------------------------


module rr_arbiter (

    input             arb_clk,      
    input             arb_rst_n,    
    input             arb_req0,  
    input             arb_req1,     
    input             arb_req2,     
    input             arb_req3,     
    output logic [1:0]  arb_gnt,
    output logic [1:0]  pointer
);

  always_ff @(posedge arb_clk or negedge arb_rst_n) begin
    if(!arb_rst_n) begin
      pointer <= 2'b00;   
      arb_gnt <= 2'b00;   
    end
    else begin
      case(pointer)
        2'b00: begin
          if(arb_req0)      arb_gnt <= 2'b00;
          else if(arb_req1) arb_gnt <= 2'b01;
          else if(arb_req2) arb_gnt <= 2'b10;
          else if(arb_req3) arb_gnt <= 2'b11;
          else              arb_gnt <= 2'b00; 
        end

        2'b01: begin
          if(arb_req1)      arb_gnt <= 2'b01;
          else if(arb_req2) arb_gnt <= 2'b10;
          else if(arb_req3) arb_gnt <= 2'b11;
          else if(arb_req0) arb_gnt <= 2'b00;
          else              arb_gnt <= 2'b00;
        end

        2'b10: begin
          if(arb_req2)      arb_gnt <= 2'b10;
          else if(arb_req3) arb_gnt <= 2'b11;
          else if(arb_req0) arb_gnt <= 2'b00;
          else if(arb_req1) arb_gnt <= 2'b01;
          else              arb_gnt <= 2'b00;
        end

        2'b11: begin
          if(arb_req3)      arb_gnt <= 2'b11;
          else if(arb_req0) arb_gnt <= 2'b00;
          else if(arb_req1) arb_gnt <= 2'b01;
          else if(arb_req2) arb_gnt <= 2'b10;
          else              arb_gnt <= 2'b00;
        end
      endcase

      pointer <= pointer + 1;
    end
  end

endmodule

//------------------------------------------------------------------------------------------------------------
//test_bench_for_assertion
//----------------------------------------------------------------------------------------------------------------------------------
module tb_rr_arbiter;

  logic arb_clk;
  logic arb_rst_n;
  logic arb_req0, arb_req1, arb_req2, arb_req3;
  logic [1:0] arb_gnt;
  logic [1:0] pointer;

  // ----------------------------------------------------------
  // DUT
  // ----------------------------------------------------------
  rr_arbiter DUT (
    .arb_clk(arb_clk),
    .arb_rst_n(arb_rst_n),
    .arb_req0(arb_req0),
    .arb_req1(arb_req1),
    .arb_req2(arb_req2),
    .arb_req3(arb_req3),
    .arb_gnt(arb_gnt),
    .pointer(pointer)
  );



  initial begin
    arb_clk = 0;
    forever #5 arb_clk = ~arb_clk;
  end

  initial begin
    arb_rst_n = 0;
    {arb_req0,arb_req1,arb_req2,arb_req3} = 4'b0000;

    #12;
    arb_rst_n = 1;

    #10 arb_req0 = 1;
    #20 arb_req1 = 1;
    #20 arb_req2 = 1;
    #20 arb_req3 = 1;
    #60 arb_req0 = 0;
    #20 arb_req1 = 0;
    #20 arb_req2 = 0;
    #20 arb_req3 = 0;

    #50 $finish;
  end

  // ----------------------------------------------------------
  // Monitor
  // ----------------------------------------------------------
  always @(posedge arb_clk) begin
    $display("T=%0t | Req0=%b,Req1=%b,Req2=%b,Req3=%b | Gnt=%b | Pointer=%b",
             $time, arb_req0,arb_req1,arb_req2,arb_req3, arb_gnt, pointer);
  end

  // ----------------------------------------------------------
  // Correct Assertions 
  // ----------------------------------------------------------

  // grant must be 0,1,2 or 3 only
   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
        arb_gnt inside {2'b00,2'b01,2'b10,2'b11})
    else $error("Invalid grant encoding");

  // Only one grant (encoded), so always true
   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
        $onehot0(1 << arb_gnt))
    else $error("Grant is not one-hot encoded!");

  // arbiter must be grant when request is high
   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
        arb_gnt==2'b00 |-> arb_req0);

   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
        arb_gnt==2'b01 |-> arb_req1);

   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
        arb_gnt==2'b10 |-> arb_req2);

   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
        arb_gnt==2'b11 |-> arb_req3);

  // Waiting time (1–4 cycles)
   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
        arb_req0 |-> ##[1:4] (arb_gnt==2'b00));

   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
        arb_req1 |-> ##[1:4] (arb_gnt==2'b01));

   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
        arb_req2 |-> ##[1:4] (arb_gnt==2'b10));

   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
        arb_req3 |-> ##[1:4] (arb_gnt==2'b11));

  // Pointer-based priority check
   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
       (pointer==2'b00 && arb_req0) |-> (arb_gnt==2'b00));

   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
       (pointer==2'b01 && arb_req1) |-> (arb_gnt==2'b01));

   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
       (pointer==2'b10 && arb_req2) |-> (arb_gnt==2'b10));

   assert property (@(posedge arb_clk) disable iff(!arb_rst_n)
       (pointer==2'b11 && arb_req3) |-> (arb_gnt==2'b11));

endmodule


